module SubBytes (
);
    
endmodule