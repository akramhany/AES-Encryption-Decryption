/*
    *
    * Module: 
    * Description:
    * ==============================================
    * Inputs:

    * Outputs:


    * Author: Akram Hany
    * Date: 10 - May - 2023 
*/

`include "slave.v"
`include "master.v"

module test_wrapper();

localparam PERIOD = 10;

localparam SIZE_128 = 8'd16;
localparam SIZE_192 = 8'd24;
localparam SIZE_256 = 8'd32;

localparam IDLE = 3'b000;
localparam SEND_ENC = 3'b001;
localparam REC_ENC = 3'b010;
localparam CHECK_ENC = 3'b011;
localparam SEND_DEC = 3'b100;
localparam REC_DEC = 3'101;
localparam CHECK_DEC = 3'b110;


/// for testing, sending and reciving data
wire [127:0] plane_text;
assign plane_text = 128'h00112233445566778899aabbccddeeff;
wire [127:0] enc_text;
assign enc_text = 128'h8ea2b7ca516745bfeafc49904b496089;
reg [127:0] test_result_send;
reg [127:0] test_result_recive;
reg [255:0] key = 256'h000102030405060708090a0b0c0d0e0f101112131415161718191a1b1c1d1e1f;


reg clk = 0;
always #(PERIOD / 2) clk = ~clk;

reg reset;
reg start;
wire buzy;
wire done;
reg [7:0] data_in;
wire [7:0] data_out;
wire cs;
wire mosi;
wire miso;
wire sclk;

wire slave_done;
reg [7:0] slave_data_in;
wire [7:0] slave_data_out;

reg start_system = 1;
reg [2:0] wrapper_state = IDLE;
reg [7:0] key_size;

master dut (
    .reset(reset),
    .clk(clk),
    .start(start),
    .buzy(buzy),
    .done(done),
    .data_in(data_in),
    .data_out(data_out),
    .cs(cs),
    .mosi(mosi),
    .miso(miso),
    .sclk(sclk)  
);

always @(posedge clk) begin

  if (reset) begin        
    wrapper_state   <= IDLE;
  end
  //TODO: put a condition to check if the start_system is 0 (make it asyncho)

end

reg [5:0] i = 0;

always @ (*)  begin

case (wrapper_state)
    
    IDLE: begin

        start = 0;
        data_in = 8'h00;
        slave_data_in = 8'h00;
        key_size = SIZE_256;
        i = key_size + 16;
        //TODO: create another reg of size 256 to store the key in it
        if (start_system && ~reset) begin
            wrapper_state = SEND_ENC;
        end
    end

    SEND_ENC: begin

        
        if (i == key_size + 16) begin
            start = 1;
            data_in = plane_text[127 -: 8];
            i = i - 1;
        end

        if (slave_done) begin
            start = 1;
            if (i > key_size)    begin
                data_in = plane_text[(i - key_size) * 8 - 1 -: 8];
                i = i - 1;
            end
            else if (i >= 0 && i < key_size)    begin
                data_in = key[(i + 1) * 8 - 1 -: 8];
                i = i - 1;
            end
            else if (i == key_size)   begin
                data_in = key_size;
                i = i - 1;
            end
            else begin
                wrapper_state = REC_ENC;
                i = 16;
            end
        end
        else begin
            start = 0;
        end
    
    end

    REC_ENC: begin

        if (slave_done) begin
            if (i > 0) begin
                start = 1;
                test_result_recive[i * 8 - 1 -: 8] = data_out;
                i = i - 1;
            end
            else    begin
                wrapper_state = CHECK_ENC;
                i = key_size + 16;
            end
        end
        else    begin
            start = 0;  //Note: think if handling start should be done in the encrypt or not
        end
    end

    CHECK_ENC: begin
        if (test_result_recive == enc_text) begin
            $display("Finallyyyyyyyyyyyyyy");
        end
        else begin
            $display("Kill me please");
        end
        start_system = 0;   //TODO: delete this statement if you want the program to run normally
        wrapper_state = IDLE;
    end

endcase
end



endmodule